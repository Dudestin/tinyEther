// Verilog netlist created by TD v4.4.433
// Wed Aug 10 04:04:58 2022

`timescale 1ns / 1ps
module sram9k  // al_ip/sram9k.v(14)
  (
  addra,
  clka,
  dia,
  rsta,
  wea,
  doa
  );

  input [9:0] addra;  // al_ip/sram9k.v(19)
  input clka;  // al_ip/sram9k.v(21)
  input [31:0] dia;  // al_ip/sram9k.v(18)
  input rsta;  // al_ip/sram9k.v(22)
  input [3:0] wea;  // al_ip/sram9k.v(20)
  output [31:0] doa;  // al_ip/sram9k.v(16)


  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0601EFE305B52500A5000C933701010101010101010101010101018100000000),
    .INIT_01(256'h83F49D2323227905F20107C47D07E417C41923220105F2980300DDF7A903A300),
    .INIT_02(256'hE770C4A4000682220107C4F4FD831123833E83638303639303A383C705F7C48A),
    .INIT_03(256'hC44913639303F447C44D13639303F407C4C913639303F4C7C4CD136393032513),
    .INIT_04(256'hC40913639303F447C40D13639303F407C48913639303F4C7C48D13639303F487),
    .INIT_05(256'h938370E750C4D123938380E7F0C4D523938390E790C4F4C7C4CD13639303F487),
    .INIT_06(256'h23C4191363C49123938340E770C49523938350E710C45123938360E7B0C45523),
    .INIT_07(256'h70E79903F4E18380E79D03F4DD8390E7A10323C4F91363C43123C4ED1363C425),
    .INIT_08(256'h03F4F58330E78903F4F18340E78D03F4ED8350E79103F4E98360E79503F4E583),
    .INIT_09(256'h8444F400A9C4AD837DB723F323A400068262D913F4FD83109183F4F98320E785),
    .INIT_0A(256'h223EA9000682223E938323B7E3C4F49C009813B700F4447103C4E707B704F4F7),
    .INIT_0B(256'h852323239323802239453E83C4C4F4B903C4F4B903C4F4B903C4F49C83232282),
    .INIT_0C(256'hC78563098484048A8304F4C4E7F084F4BA8303AA3E93B303842D232383F48587),
    .INIT_0D(256'hE393032304E7F704BA038304E784C4F485838785E39303234444E947853E8A83),
    .INIT_0E(256'h91B723B7220121628113E7F0C4F485838513459183C7856393831383C4C49923),
    .INIT_0F(256'h8785478547850785010785478587850785C7854785C7854785E33E3D13012380),
    .INIT_10(256'h308262014785C785478507850785C785878587858785878587858785C7854785),
    .INIT_11(256'h74547350007320742A594546202E0A742A4F45462000656D6952303E00633834),
    .INIT_12(256'h7C20205F5F5F205F207C205F205F5F5F5F5F200A5F20205F20205F5F202E6E6F),
    .INIT_13(256'h203A746E63530A203A6D6C547C5F5F205F5F5F5F20200A7C297C5F5F5F205F20),
    .INIT_14(256'h3520644F6C2068773420652061206877332000656943536532200A6846536531),
    .INIT_15(256'h00616E636969753920646420756E656F37206452642068773620644F64206877),
    .INIT_16(256'h00000000000000000A556365207420207253207365754D200A6620206D653020),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_1024x32_sub_000000_000 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia({open_n69,dia[7:0]}),
    .rsta(rsta),
    .wea(wea[0]),
    .doa({open_n83,doa[7:0]}));
  // address_offset=0;data_offset=8;depth=1024;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hCEA0004D0000B000B000C105054F4E4D4C4B4A49484746454443424000000000),
    .INIT_01(256'h27FE472C2ED47161400000FE3700FE00FEA826CC116140C34702370047470710),
    .INIT_02(256'h003EFEFE10CE805400FAFEFE1727A02C2785475B272718074705C7876700FD07),
    .INIT_03(256'hFE3505FC0727FED4FE3505FC0727FECEFE3505FC0727FEC7FE3505FC07273785),
    .INIT_04(256'hFE3505FC0727FEEDFE3505FC0727FEE7FE3505FC0727FEE0FE3505FC0727FEDA),
    .INIT_05(256'h8727030004FEA8268727030004FEA8268727030005FEFEF9FE3305FB0727FEF3),
    .INIT_06(256'h26FE3305FBFEA8268727030002FEA8268727030003FEA8268727030003FEA826),
    .INIT_07(256'h03004727FE172703004727FE17270300472726FE3105FAFEA826FE3105FBFEA8),
    .INIT_08(256'h27FE172703004727FE172703004727FE172703004727FE172703004727FE1727),
    .INIT_09(256'hFEFEFEC0A8FDC3275707242726FC18D680443605FE172703CB27FE1727030047),
    .INIT_0A(256'h44853708C6805485F727A00701FEFE4302C3470703FEFE3625FD02B000FEFE40),
    .INIT_0B(256'h6726282A072C00DC71618527FEFDFE8F27FEFE8F27FEFE8F27FEFE43272ED680),
    .INIT_0C(256'h8A67813FFC43FD0727FEFCFEFC03FEFE9727278785070427FEA0242427FE4789),
    .INIT_0D(256'hDC072720FE000FFE972727FEF4FDFEFE07278C67F8072722FDFEA08C67850727),
    .INIT_0E(256'h0707A007CC1161543A85FA07FDFC07273A853A45278C6700F727F7C7FCFDA02E),
    .INIT_0F(256'h9E678C678C679E67459D678C679A6798679567936790678C6719873385002606),
    .INIT_10(256'h318044008C67B467B367B267B067AD67AB67A967A767A567A367A1679F678C67),
    .INIT_11(256'h6F452072006570202A5444412A0000202A5244412A0073656E75303D00643935),
    .INIT_12(256'h0A5C2F5F205F7C297C0A5F20205F5F5F29207C005F20205F2020205F200A756E),
    .INIT_13(256'h200A69207465004B206F206F0A5F2F5C5F5F5F7C207C005F20205F297C7C5F7C),
    .INIT_14(256'h5D206520204420695D200A6D756420695D200067676F50615D2000206C50615D),
    .INIT_15(256'h00726320736D6E5D206520726F7420675D206520205120695D20652020512069),
    .INIT_16(256'h00000000000000000041685D20657353695D20746D6E5D2000696361616E5D20),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_1024x32_sub_000000_008 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia({open_n115,dia[15:8]}),
    .rsta(rsta),
    .wea(wea[1]),
    .doa({open_n129,doa[15:8]}));
  // address_offset=0;data_offset=16;depth=1024;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h220140B511236393971317F00081818181818181818181818181818100000000),
    .INIT_01(256'hC4A123B4A40006826201F583833E83231383A40006826201F4A1B73563F4F4AA),
    .INIT_02(256'h8563930323220145B201E38323C401F4C481B4F784C4F700B4F407BA13BDB303),
    .INIT_03(256'h938360E770C4C123938370E7B0C4C523938380E7F0C40123938390E730C40507),
    .INIT_04(256'h938320E770C48123938330E7B0C48523938340E7F0C44123938350E730C44523),
    .INIT_05(256'hA7C45113639303F407C45513639303F467C4D11363930323938310E730C40523),
    .INIT_06(256'hF4898330E7F503F487C41513639303F4E7C49113639303F447C49513639303F4),
    .INIT_07(256'hB51363C4E123C4611363C4D523C4551363C4F4D98310E7A503F4B18320E7CD03),
    .INIT_08(256'hC43523C4311363C4A123C4251363C49523C4911363C44123C4851363C47523C4),
    .INIT_09(256'hB3830323F3C903C49800F400F4FD23227905F2002123C4E113C40523C4C51363),
    .INIT_0A(256'h41B2AA01224145B2F7C40700F7FD0323A1B7F70098B72383C481836393B70323),
    .INIT_0B(256'h130404F400F49526068232C498038323C4968323C4C58323C4B68323C4A40079),
    .INIT_0C(256'h3D13F4AA3E93BA0344A9232383E393032344849C9184F7048A8304F4C465236D),
    .INIT_0D(256'hE7F004F48583231303C4040D23E3830323C4DD13E7F044F4BA83032913A99144),
    .INIT_0E(256'h13000700000682D2F24785E3930323C40547853EC44913F7F7C4F707BA038304),
    .INIT_0F(256'h7D135D137D13D91361C913E913CD13ED13CD13ED1309132913F7B5AA07850498),
    .INIT_10(256'h320005F23D139913B9139913B9139D13BD139D13BD1359137913591379135D13),
    .INIT_11(256'h2052456500646100204520492A000000204420492A00746D676E003100656136),
    .INIT_12(256'h007C20205C2F2F2020005F205F5F2F20205C20005F20205F202020205F006574),
    .INIT_13(256'h20006F61206C006900726D74005F205F5F2F5C5C205F005F7C28292020202F20),
    .INIT_14(256'h20200A6D497574742020006F6C65747420200073206E49642020004961496420),
    .INIT_15(256'h006B686274702020200A6D657569636720200A6D4475747420200A6D49757474),
    .INIT_16(256'h000000000000000000526F20200A74506E20200A7420202000676F6C72632020),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_1024x32_sub_000000_016 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia({open_n161,dia[23:16]}),
    .rsta(rsta),
    .wea(wea[2]),
    .doa({open_n175,doa[23:16]}));
  // address_offset=0;data_offset=24;depth=1024;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hCC116FFE05205785150515FF034F4E4D4C4B4A49484746454443424100000000),
    .INIT_01(256'hFEA826FCFC18D6804400F3C72785C7268727FE10CE804400FE07074514FEFE87),
    .INIT_02(256'h67F7072726CC11615000D32726FE00FCFE37FE00FDFE0003FEFE0097078B5727),
    .INIT_03(256'h8727030025FEA026872703002BFEA0268727030031FEA2268727030038FEAE89),
    .INIT_04(256'h872703000CFEA0268727030012FEA0268727030018FEA026872703001FFEA026),
    .INIT_05(256'hFBFE3305FC0727FEFBFE3305FC0727FEFAFE3305FC0727268727030006FEA026),
    .INIT_06(256'hFE172703004727FEFDFE3305FC0727FEFCFE3305FC0727FEFCFE3305FC0727FE),
    .INIT_07(256'h3905FBFEA026FE3905FBFEA026FE3905FBFEFE172703004727FE172703004727),
    .INIT_08(256'hFEA826FE3105FBFEA826FE3105FBFEA826FE3105FBFEA826FE3105FBFEA026FE),
    .INIT_09(256'h07272722273625FDC303FEC0FE572ED471614003A026FE3E05FEA026FE3E05FB),
    .INIT_0A(256'h01408745C41161500FFE0003FA5727260707FF0343072427FDC727F487272720),
    .INIT_0B(256'h85FCFCFC10FC47DADE8054FEC3272726FE072726FE832726FE072726FDFC1871),
    .INIT_0C(256'h3485028785079727FEA0222427F8072724FDFEC03FFC00FD0727FEFCFEA82634),
    .INIT_0D(256'hFC07FEFE0727807727FCFEA020D1272726FE3A85FA03FEFE9727273C853C45FE),
    .INIT_0E(256'h0702000310CE8054508E67DA07272EFDA08C6785FD3285020FFD0F00972727FC),
    .INIT_0F(256'h30853885388530853238853885308530853885388532853285FE47878F67FEC3),
    .INIT_10(256'h3300614038853085308538853885308530853885388530853085388538853085),
    .INIT_11(256'h63204E73000A7300612A424C2A000000612A574C2A002074206E003000666237),
    .INIT_12(256'h00205F5C5F20207C7C005F2F5F7C205F5F2820005F2020205F2020205F002E69),
    .INIT_13(256'h5B006E636165004200796561005F5C5F2F5F5F5F7C7C005F205F207C28287C20),
    .INIT_14(256'h535B006F2F616F63535B006474666F63535B000A52662020525B004473202052),
    .INIT_15(256'h000A6D65696C73525B006F61736E6F6C545B006F44616F63535B006F2F616F63),
    .INIT_16(256'h0000000000000000005420455B00614974505B00654D525B00736E6C6B68425B),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_1024x32_sub_000000_024 (
    .addra({addra,3'b111}),
    .clka(clka),
    .dia({open_n207,dia[31:24]}),
    .rsta(rsta),
    .wea(wea[3]),
    .doa({open_n221,doa[31:24]}));

endmodule 

